sleebarr@sleebarr-Inspiron-3420.11067:1509028106